* A voltage divider circuit

* Sinusoidal input
V1 1 0 SIN (0 1 1k)

* Resistors
R1 1 2 1k
R2 2 0 1k

* Transient Simulation
.tran 1u 1m

.end
